`ifndef _DEFINES_H_
`define _DEFINES_H_

// Parameters
// `define {name} {value}


// Instruction Memory

`define IMEM_ADDR_WIDTH 32
`define IMEM_DATA_WIDTH 32
`define IMEM_WIDTH 8
`define IMEM_DEPTH 256

`endif